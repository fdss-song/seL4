arch x86_64

objects {
buf2_frame_cap = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 102400}])
cnode_threads = cnode (4 bits)
frame_threads_0000 = frame (4k, fill: [{0 548 CDL_FrameFill_FileData "threads" 0}])
frame_threads_0001 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 4096}])
frame_threads_0002 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 8192}])
frame_threads_0003 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 12288}])
frame_threads_0004 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 16384}])
frame_threads_0005 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 20480}])
frame_threads_0006 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 24576}])
frame_threads_0007 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 28672}])
frame_threads_0008 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 32768}])
frame_threads_0009 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 36864}])
frame_threads_0010 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 40960}])
frame_threads_0011 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 45056}])
frame_threads_0012 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 49152}])
frame_threads_0013 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 53248}])
frame_threads_0014 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 57344}])
frame_threads_0015 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 61440}])
frame_threads_0016 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 65536}])
frame_threads_0017 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 69632}])
frame_threads_0018 = frame (4k, fill: [{0 582 CDL_FrameFill_FileData "threads" 73728}])
frame_threads_0019 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 77824}])
frame_threads_0020 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 81920}])
frame_threads_0021 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 86016}])
frame_threads_0022 = frame (4k, fill: [{0 2672 CDL_FrameFill_FileData "threads" 90112}])
frame_threads_0023 = frame (4k, fill: [{4040 56 CDL_FrameFill_FileData "threads" 94152}])
frame_threads_0024 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 94208}])
frame_threads_0025 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 98304}])
frame_threads_0028 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 110592}])
frame_threads_0029 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 114688}])
frame_threads_0030 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 118784}])
frame_threads_0031 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 122880}])
frame_threads_0032 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 126976}])
frame_threads_0033 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 131072}])
frame_threads_0034 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 135168}])
frame_threads_0035 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 139264}])
frame_threads_0036 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 143360}])
frame_threads_0037 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 147456}])
frame_threads_0038 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 151552}])
frame_threads_0039 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 155648}])
frame_threads_0040 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 159744}])
frame_threads_0041 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 163840}])
frame_threads_0042 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 167936}])
frame_threads_0043 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 172032}])
frame_threads_0061 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "threads" 245760}])
frame_threads_0062 = frame (4k, fill: [])
frame_threads_0063 = frame (4k, fill: [])
frame_threads_0064 = frame (4k, fill: [])
frame_threads_0065 = frame (4k, fill: [])
frame_threads_0066 = frame (4k, fill: [])
frame_threads_0067 = frame (4k, fill: [])
frame_threads_0068 = frame (4k, fill: [])
frame_threads_0069 = frame (4k, fill: [])
frame_threads_0070 = frame (4k, fill: [])
frame_threads_0071 = frame (4k, fill: [])
frame_threads_0072 = frame (4k, fill: [])
frame_threads_0073 = frame (4k, fill: [])
frame_threads_0074 = frame (4k, fill: [])
frame_threads_0075 = frame (4k, fill: [])
frame_threads_0076 = frame (4k, fill: [])
frame_threads_0077 = frame (4k, fill: [])
frame_threads_0078 = frame (4k, fill: [])
frame_threads_0079 = frame (4k, fill: [])
frame_threads_0080 = frame (4k, fill: [])
frame_threads_0081 = frame (4k, fill: [])
frame_threads_0082 = frame (4k, fill: [])
frame_threads_0083 = frame (4k, fill: [])
frame_threads_0084 = frame (4k, fill: [])
frame_threads_0085 = frame (4k, fill: [])
frame_threads_0086 = frame (4k, fill: [])
frame_threads_0087 = frame (4k, fill: [])
frame_threads_0088 = frame (4k, fill: [])
frame_threads_0089 = frame (4k, fill: [])
frame_threads_0090 = frame (4k, fill: [])
frame_threads_0091 = frame (4k, fill: [])
frame_threads_0092 = frame (4k, fill: [])
frame_threads_0093 = frame (4k, fill: [])
frame_threads_0094 = frame (4k, fill: [])
frame_threads_0095 = frame (4k, fill: [])
frame_threads_0096 = frame (4k, fill: [])
frame_threads_0097 = frame (4k, fill: [])
frame_threads_0098 = frame (4k, fill: [])
frame_threads_0099 = frame (4k, fill: [])
frame_threads_0100 = frame (4k, fill: [])
frame_threads_0101 = frame (4k, fill: [])
frame_threads_0102 = frame (4k, fill: [])
frame_threads_0103 = frame (4k, fill: [])
frame_threads_0104 = frame (4k, fill: [])
frame_threads_0105 = frame (4k, fill: [])
frame_threads_0106 = frame (4k, fill: [])
frame_threads_0107 = frame (4k, fill: [])
frame_threads_0108 = frame (4k, fill: [])
frame_threads_0109 = frame (4k, fill: [])
frame_threads_0110 = frame (4k, fill: [])
frame_threads_0111 = frame (4k, fill: [])
frame_threads_0112 = frame (4k, fill: [])
frame_threads_0113 = frame (4k, fill: [])
frame_threads_0114 = frame (4k, fill: [])
frame_threads_0115 = frame (4k, fill: [])
frame_threads_0116 = frame (4k, fill: [])
frame_threads_0117 = frame (4k, fill: [])
frame_threads_0118 = frame (4k, fill: [])
frame_threads_0119 = frame (4k, fill: [])
frame_threads_0120 = frame (4k, fill: [])
frame_threads_0121 = frame (4k, fill: [])
frame_threads_0122 = frame (4k, fill: [])
frame_threads_0123 = frame (4k, fill: [])
frame_threads_0124 = frame (4k, fill: [])
frame_threads_0125 = frame (4k, fill: [])
frame_threads_0126 = frame (4k, fill: [])
frame_threads_0127 = frame (4k, fill: [])
frame_threads_0128 = frame (4k, fill: [])
frame_threads_0129 = frame (4k, fill: [])
frame_threads_0130 = frame (4k, fill: [])
frame_threads_0131 = frame (4k, fill: [])
frame_threads_0132 = frame (4k, fill: [])
frame_threads_0133 = frame (4k, fill: [])
frame_threads_0134 = frame (4k, fill: [])
frame_threads_0135 = frame (4k, fill: [])
frame_threads_0136 = frame (4k, fill: [])
frame_threads_0137 = frame (4k, fill: [])
frame_threads_0138 = frame (4k, fill: [])
frame_threads_0139 = frame (4k, fill: [])
frame_threads_0140 = frame (4k, fill: [])
frame_threads_0141 = frame (4k, fill: [])
frame_threads_0142 = frame (4k, fill: [])
frame_threads_0143 = frame (4k, fill: [])
frame_threads_0144 = frame (4k, fill: [])
frame_threads_0145 = frame (4k, fill: [])
frame_threads_0146 = frame (4k, fill: [])
frame_threads_0147 = frame (4k, fill: [])
frame_threads_0148 = frame (4k, fill: [])
frame_threads_0149 = frame (4k, fill: [])
frame_threads_0150 = frame (4k, fill: [])
frame_threads_0151 = frame (4k, fill: [])
frame_threads_0152 = frame (4k, fill: [])
frame_threads_0153 = frame (4k, fill: [])
frame_threads_0154 = frame (4k, fill: [])
frame_threads_0155 = frame (4k, fill: [])
frame_threads_0156 = frame (4k, fill: [])
frame_threads_0157 = frame (4k, fill: [])
frame_threads_0158 = frame (4k, fill: [])
frame_threads_0159 = frame (4k, fill: [])
frame_threads_0160 = frame (4k, fill: [])
frame_threads_0161 = frame (4k, fill: [])
frame_threads_0162 = frame (4k, fill: [])
frame_threads_0163 = frame (4k, fill: [])
frame_threads_0164 = frame (4k, fill: [])
frame_threads_0165 = frame (4k, fill: [])
frame_threads_0166 = frame (4k, fill: [])
frame_threads_0167 = frame (4k, fill: [])
frame_threads_0168 = frame (4k, fill: [])
frame_threads_0169 = frame (4k, fill: [])
frame_threads_0170 = frame (4k, fill: [])
frame_threads_0171 = frame (4k, fill: [])
frame_threads_0172 = frame (4k, fill: [])
frame_threads_0173 = frame (4k, fill: [])
frame_threads_0174 = frame (4k, fill: [])
frame_threads_0175 = frame (4k, fill: [])
frame_threads_0176 = frame (4k, fill: [])
frame_threads_0177 = frame (4k, fill: [])
frame_threads_0178 = frame (4k, fill: [])
frame_threads_0179 = frame (4k, fill: [])
frame_threads_0180 = frame (4k, fill: [])
frame_threads_0181 = frame (4k, fill: [])
frame_threads_0182 = frame (4k, fill: [])
frame_threads_0183 = frame (4k, fill: [])
frame_threads_0184 = frame (4k, fill: [])
frame_threads_0185 = frame (4k, fill: [])
frame_threads_0186 = frame (4k, fill: [])
frame_threads_0187 = frame (4k, fill: [])
frame_threads_0188 = frame (4k, fill: [])
frame_threads_0189 = frame (4k, fill: [])
frame_threads_0190 = frame (4k, fill: [])
frame_threads_0191 = frame (4k, fill: [])
frame_threads_0192 = frame (4k, fill: [])
frame_threads_0193 = frame (4k, fill: [])
frame_threads_0194 = frame (4k, fill: [])
frame_threads_0195 = frame (4k, fill: [])
frame_threads_0196 = frame (4k, fill: [])
frame_threads_0197 = frame (4k, fill: [])
frame_threads_0198 = frame (4k, fill: [])
frame_threads_0199 = frame (4k, fill: [])
frame_threads_0200 = frame (4k, fill: [])
frame_threads_0201 = frame (4k, fill: [])
frame_threads_0202 = frame (4k, fill: [])
frame_threads_0203 = frame (4k, fill: [])
frame_threads_0204 = frame (4k, fill: [])
frame_threads_0205 = frame (4k, fill: [])
frame_threads_0206 = frame (4k, fill: [])
frame_threads_0207 = frame (4k, fill: [])
frame_threads_0208 = frame (4k, fill: [])
frame_threads_0209 = frame (4k, fill: [])
frame_threads_0210 = frame (4k, fill: [])
frame_threads_0211 = frame (4k, fill: [])
frame_threads_0212 = frame (4k, fill: [])
frame_threads_0213 = frame (4k, fill: [])
frame_threads_0214 = frame (4k, fill: [])
frame_threads_0215 = frame (4k, fill: [])
frame_threads_0216 = frame (4k, fill: [])
frame_threads_0217 = frame (4k, fill: [])
frame_threads_0218 = frame (4k, fill: [])
frame_threads_0219 = frame (4k, fill: [])
frame_threads_0220 = frame (4k, fill: [])
frame_threads_0221 = frame (4k, fill: [])
frame_threads_0222 = frame (4k, fill: [])
frame_threads_0223 = frame (4k, fill: [])
frame_threads_0224 = frame (4k, fill: [])
frame_threads_0225 = frame (4k, fill: [])
frame_threads_0226 = frame (4k, fill: [])
frame_threads_0227 = frame (4k, fill: [])
frame_threads_0228 = frame (4k, fill: [])
frame_threads_0229 = frame (4k, fill: [])
frame_threads_0230 = frame (4k, fill: [])
frame_threads_0231 = frame (4k, fill: [])
frame_threads_0232 = frame (4k, fill: [])
frame_threads_0233 = frame (4k, fill: [])
frame_threads_0234 = frame (4k, fill: [])
frame_threads_0235 = frame (4k, fill: [])
frame_threads_0236 = frame (4k, fill: [])
frame_threads_0237 = frame (4k, fill: [])
frame_threads_0238 = frame (4k, fill: [])
frame_threads_0239 = frame (4k, fill: [])
frame_threads_0240 = frame (4k, fill: [])
frame_threads_0241 = frame (4k, fill: [])
frame_threads_0242 = frame (4k, fill: [])
frame_threads_0243 = frame (4k, fill: [])
frame_threads_0244 = frame (4k, fill: [])
frame_threads_0245 = frame (4k, fill: [])
frame_threads_0246 = frame (4k, fill: [])
frame_threads_0247 = frame (4k, fill: [])
frame_threads_0248 = frame (4k, fill: [])
frame_threads_0249 = frame (4k, fill: [])
frame_threads_0250 = frame (4k, fill: [])
frame_threads_0251 = frame (4k, fill: [])
frame_threads_0252 = frame (4k, fill: [])
frame_threads_0253 = frame (4k, fill: [])
frame_threads_0254 = frame (4k, fill: [])
frame_threads_0255 = frame (4k, fill: [])
frame_threads_0256 = frame (4k, fill: [])
frame_threads_0257 = frame (4k, fill: [])
frame_threads_0258 = frame (4k, fill: [])
frame_threads_0259 = frame (4k, fill: [])
frame_threads_0260 = frame (4k, fill: [])
frame_threads_0261 = frame (4k, fill: [])
frame_threads_0262 = frame (4k, fill: [])
frame_threads_0263 = frame (4k, fill: [])
frame_threads_0264 = frame (4k, fill: [])
frame_threads_0265 = frame (4k, fill: [])
frame_threads_0266 = frame (4k, fill: [])
frame_threads_0267 = frame (4k, fill: [])
frame_threads_0268 = frame (4k, fill: [])
frame_threads_0269 = frame (4k, fill: [])
frame_threads_0270 = frame (4k, fill: [])
frame_threads_0271 = frame (4k, fill: [])
frame_threads_0272 = frame (4k, fill: [])
frame_threads_0273 = frame (4k, fill: [])
frame_threads_0274 = frame (4k, fill: [])
frame_threads_0275 = frame (4k, fill: [])
frame_threads_0276 = frame (4k, fill: [])
frame_threads_0277 = frame (4k, fill: [])
frame_threads_0278 = frame (4k, fill: [])
frame_threads_0279 = frame (4k, fill: [])
frame_threads_0280 = frame (4k, fill: [])
frame_threads_0281 = frame (4k, fill: [])
frame_threads_0282 = frame (4k, fill: [])
frame_threads_0283 = frame (4k, fill: [])
frame_threads_0284 = frame (4k, fill: [])
frame_threads_0285 = frame (4k, fill: [])
frame_threads_0286 = frame (4k, fill: [])
frame_threads_0287 = frame (4k, fill: [])
frame_threads_0288 = frame (4k, fill: [])
frame_threads_0289 = frame (4k, fill: [])
frame_threads_0290 = frame (4k, fill: [])
frame_threads_0291 = frame (4k, fill: [])
frame_threads_0292 = frame (4k, fill: [])
frame_threads_0293 = frame (4k, fill: [])
frame_threads_0294 = frame (4k, fill: [])
frame_threads_0295 = frame (4k, fill: [])
frame_threads_0296 = frame (4k, fill: [])
frame_threads_0297 = frame (4k, fill: [])
frame_threads_0298 = frame (4k, fill: [])
frame_threads_0299 = frame (4k, fill: [])
frame_threads_0300 = frame (4k, fill: [])
frame_threads_0301 = frame (4k, fill: [])
frame_threads_0302 = frame (4k, fill: [])
frame_threads_0303 = frame (4k, fill: [])
frame_threads_0304 = frame (4k, fill: [])
frame_threads_0305 = frame (4k, fill: [])
frame_threads_0306 = frame (4k, fill: [])
frame_threads_0307 = frame (4k, fill: [])
frame_threads_0308 = frame (4k, fill: [])
frame_threads_0309 = frame (4k, fill: [])
frame_threads_0310 = frame (4k, fill: [])
frame_threads_0311 = frame (4k, fill: [])
frame_threads_0312 = frame (4k, fill: [])
frame_threads_0313 = frame (4k, fill: [])
frame_threads_0314 = frame (4k, fill: [])
frame_threads_0315 = frame (4k, fill: [])
frame_threads_0316 = frame (4k, fill: [])
frame_threads_0317 = frame (4k, fill: [])
frame_threads_0318 = frame (4k, fill: [])
frame_threads_0319 = frame (4k, fill: [])
frame_threads_0320 = frame (4k, fill: [])
frame_threads_0321 = frame (4k, fill: [])
frame_threads_0322 = frame (4k, fill: [])
frame_threads_0323 = frame (4k, fill: [])
frame_threads_0324 = frame (4k, fill: [])
ipc_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 241664}])
pd_threads_0001 = pd
pdpt_threads_0000 = pdpt
pt_threads_0002 = pt
stack_0_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 176128}])
stack_10_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 217088}])
stack_11_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 221184}])
stack_12_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 225280}])
stack_13_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 229376}])
stack_14_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 233472}])
stack_15_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 237568}])
stack_1_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 180224}])
stack_2_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 184320}])
stack_3_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 188416}])
stack_4_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 192512}])
stack_5_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 196608}])
stack_6_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 200704}])
stack_7_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 204800}])
stack_8_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 208896}])
stack_9_threads_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 212992}])
tcb_ipc_frame = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "threads" 106496}])
tcb_threads = tcb (addr: 0x43c000,ip: 0x401034,sp: 0x42d000,prio: 254,max_prio: 254,affinity: 0,init: [0, 0, 0, 0, 2, 4292672, 1, 0, 0, 32, 4212419, 0, 0])
tcb_untyped = ut (11 bits) {  }
vspace_threads = pml4
}

caps {
cnode_threads {
0x1: cnode_threads (guard: 0, guard_size: 60)
0x2: vspace_threads
0x3: tcb_threads
0x4: tcb_untyped
0x5: buf2_frame_cap (RWX)
0x7: tcb_ipc_frame (RWX)
0x8: tcb_threads
}
pd_threads_0001 {
0x2: pt_threads_0002
}
pdpt_threads_0000 {
0x0: pd_threads_0001
}
pt_threads_0002 {
0x0: frame_threads_0000 (R)
0x1: frame_threads_0001 (RX)
0x2: frame_threads_0002 (RX)
0x3: frame_threads_0003 (RX)
0x4: frame_threads_0004 (RX)
0x5: frame_threads_0005 (RX)
0x6: frame_threads_0006 (RX)
0x7: frame_threads_0007 (RX)
0x8: frame_threads_0008 (RX)
0x9: frame_threads_0009 (RX)
0xa: frame_threads_0010 (RX)
0xb: frame_threads_0011 (RX)
0xc: frame_threads_0012 (RX)
0xd: frame_threads_0013 (RX)
0xe: frame_threads_0014 (RX)
0xf: frame_threads_0015 (RX)
0x10: frame_threads_0016 (RX)
0x11: frame_threads_0017 (RX)
0x12: frame_threads_0018 (RX)
0x13: frame_threads_0019 (R)
0x14: frame_threads_0020 (R)
0x15: frame_threads_0021 (R)
0x16: frame_threads_0022 (R)
0x17: frame_threads_0023 (RW)
0x18: frame_threads_0024 (RW)
0x19: frame_threads_0025 (RW)
0x1a: buf2_frame_cap (RWX)
0x1b: tcb_ipc_frame (RWX)
0x1c: frame_threads_0028 (RW)
0x1d: frame_threads_0029 (RW)
0x1e: frame_threads_0030 (RW)
0x1f: frame_threads_0031 (RW)
0x20: frame_threads_0032 (RW)
0x21: frame_threads_0033 (RW)
0x22: frame_threads_0034 (RW)
0x23: frame_threads_0035 (RW)
0x24: frame_threads_0036 (RW)
0x25: frame_threads_0037 (RW)
0x26: frame_threads_0038 (RW)
0x27: frame_threads_0039 (RW)
0x28: frame_threads_0040 (RW)
0x29: frame_threads_0041 (RW)
0x2a: frame_threads_0042 (RW)
0x2b: frame_threads_0043 (RW)
0x2c: stack_0_threads_obj (RW)
0x2d: stack_1_threads_obj (RW)
0x2e: stack_2_threads_obj (RW)
0x2f: stack_3_threads_obj (RW)
0x30: stack_4_threads_obj (RW)
0x31: stack_5_threads_obj (RW)
0x32: stack_6_threads_obj (RW)
0x33: stack_7_threads_obj (RW)
0x34: stack_8_threads_obj (RW)
0x35: stack_9_threads_obj (RW)
0x36: stack_10_threads_obj (RW)
0x37: stack_11_threads_obj (RW)
0x38: stack_12_threads_obj (RW)
0x39: stack_13_threads_obj (RW)
0x3a: stack_14_threads_obj (RW)
0x3b: stack_15_threads_obj (RW)
0x3c: ipc_threads_obj (RW)
0x3d: frame_threads_0061 (RW)
0x3e: frame_threads_0062 (RW)
0x3f: frame_threads_0063 (RW)
0x40: frame_threads_0064 (RW)
0x41: frame_threads_0065 (RW)
0x42: frame_threads_0066 (RW)
0x43: frame_threads_0067 (RW)
0x44: frame_threads_0068 (RW)
0x45: frame_threads_0069 (RW)
0x46: frame_threads_0070 (RW)
0x47: frame_threads_0071 (RW)
0x48: frame_threads_0072 (RW)
0x49: frame_threads_0073 (RW)
0x4a: frame_threads_0074 (RW)
0x4b: frame_threads_0075 (RW)
0x4c: frame_threads_0076 (RW)
0x4d: frame_threads_0077 (RW)
0x4e: frame_threads_0078 (RW)
0x4f: frame_threads_0079 (RW)
0x50: frame_threads_0080 (RW)
0x51: frame_threads_0081 (RW)
0x52: frame_threads_0082 (RW)
0x53: frame_threads_0083 (RW)
0x54: frame_threads_0084 (RW)
0x55: frame_threads_0085 (RW)
0x56: frame_threads_0086 (RW)
0x57: frame_threads_0087 (RW)
0x58: frame_threads_0088 (RW)
0x59: frame_threads_0089 (RW)
0x5a: frame_threads_0090 (RW)
0x5b: frame_threads_0091 (RW)
0x5c: frame_threads_0092 (RW)
0x5d: frame_threads_0093 (RW)
0x5e: frame_threads_0094 (RW)
0x5f: frame_threads_0095 (RW)
0x60: frame_threads_0096 (RW)
0x61: frame_threads_0097 (RW)
0x62: frame_threads_0098 (RW)
0x63: frame_threads_0099 (RW)
0x64: frame_threads_0100 (RW)
0x65: frame_threads_0101 (RW)
0x66: frame_threads_0102 (RW)
0x67: frame_threads_0103 (RW)
0x68: frame_threads_0104 (RW)
0x69: frame_threads_0105 (RW)
0x6a: frame_threads_0106 (RW)
0x6b: frame_threads_0107 (RW)
0x6c: frame_threads_0108 (RW)
0x6d: frame_threads_0109 (RW)
0x6e: frame_threads_0110 (RW)
0x6f: frame_threads_0111 (RW)
0x70: frame_threads_0112 (RW)
0x71: frame_threads_0113 (RW)
0x72: frame_threads_0114 (RW)
0x73: frame_threads_0115 (RW)
0x74: frame_threads_0116 (RW)
0x75: frame_threads_0117 (RW)
0x76: frame_threads_0118 (RW)
0x77: frame_threads_0119 (RW)
0x78: frame_threads_0120 (RW)
0x79: frame_threads_0121 (RW)
0x7a: frame_threads_0122 (RW)
0x7b: frame_threads_0123 (RW)
0x7c: frame_threads_0124 (RW)
0x7d: frame_threads_0125 (RW)
0x7e: frame_threads_0126 (RW)
0x7f: frame_threads_0127 (RW)
0x80: frame_threads_0128 (RW)
0x81: frame_threads_0129 (RW)
0x82: frame_threads_0130 (RW)
0x83: frame_threads_0131 (RW)
0x84: frame_threads_0132 (RW)
0x85: frame_threads_0133 (RW)
0x86: frame_threads_0134 (RW)
0x87: frame_threads_0135 (RW)
0x88: frame_threads_0136 (RW)
0x89: frame_threads_0137 (RW)
0x8a: frame_threads_0138 (RW)
0x8b: frame_threads_0139 (RW)
0x8c: frame_threads_0140 (RW)
0x8d: frame_threads_0141 (RW)
0x8e: frame_threads_0142 (RW)
0x8f: frame_threads_0143 (RW)
0x90: frame_threads_0144 (RW)
0x91: frame_threads_0145 (RW)
0x92: frame_threads_0146 (RW)
0x93: frame_threads_0147 (RW)
0x94: frame_threads_0148 (RW)
0x95: frame_threads_0149 (RW)
0x96: frame_threads_0150 (RW)
0x97: frame_threads_0151 (RW)
0x98: frame_threads_0152 (RW)
0x99: frame_threads_0153 (RW)
0x9a: frame_threads_0154 (RW)
0x9b: frame_threads_0155 (RW)
0x9c: frame_threads_0156 (RW)
0x9d: frame_threads_0157 (RW)
0x9e: frame_threads_0158 (RW)
0x9f: frame_threads_0159 (RW)
0xa0: frame_threads_0160 (RW)
0xa1: frame_threads_0161 (RW)
0xa2: frame_threads_0162 (RW)
0xa3: frame_threads_0163 (RW)
0xa4: frame_threads_0164 (RW)
0xa5: frame_threads_0165 (RW)
0xa6: frame_threads_0166 (RW)
0xa7: frame_threads_0167 (RW)
0xa8: frame_threads_0168 (RW)
0xa9: frame_threads_0169 (RW)
0xaa: frame_threads_0170 (RW)
0xab: frame_threads_0171 (RW)
0xac: frame_threads_0172 (RW)
0xad: frame_threads_0173 (RW)
0xae: frame_threads_0174 (RW)
0xaf: frame_threads_0175 (RW)
0xb0: frame_threads_0176 (RW)
0xb1: frame_threads_0177 (RW)
0xb2: frame_threads_0178 (RW)
0xb3: frame_threads_0179 (RW)
0xb4: frame_threads_0180 (RW)
0xb5: frame_threads_0181 (RW)
0xb6: frame_threads_0182 (RW)
0xb7: frame_threads_0183 (RW)
0xb8: frame_threads_0184 (RW)
0xb9: frame_threads_0185 (RW)
0xba: frame_threads_0186 (RW)
0xbb: frame_threads_0187 (RW)
0xbc: frame_threads_0188 (RW)
0xbd: frame_threads_0189 (RW)
0xbe: frame_threads_0190 (RW)
0xbf: frame_threads_0191 (RW)
0xc0: frame_threads_0192 (RW)
0xc1: frame_threads_0193 (RW)
0xc2: frame_threads_0194 (RW)
0xc3: frame_threads_0195 (RW)
0xc4: frame_threads_0196 (RW)
0xc5: frame_threads_0197 (RW)
0xc6: frame_threads_0198 (RW)
0xc7: frame_threads_0199 (RW)
0xc8: frame_threads_0200 (RW)
0xc9: frame_threads_0201 (RW)
0xca: frame_threads_0202 (RW)
0xcb: frame_threads_0203 (RW)
0xcc: frame_threads_0204 (RW)
0xcd: frame_threads_0205 (RW)
0xce: frame_threads_0206 (RW)
0xcf: frame_threads_0207 (RW)
0xd0: frame_threads_0208 (RW)
0xd1: frame_threads_0209 (RW)
0xd2: frame_threads_0210 (RW)
0xd3: frame_threads_0211 (RW)
0xd4: frame_threads_0212 (RW)
0xd5: frame_threads_0213 (RW)
0xd6: frame_threads_0214 (RW)
0xd7: frame_threads_0215 (RW)
0xd8: frame_threads_0216 (RW)
0xd9: frame_threads_0217 (RW)
0xda: frame_threads_0218 (RW)
0xdb: frame_threads_0219 (RW)
0xdc: frame_threads_0220 (RW)
0xdd: frame_threads_0221 (RW)
0xde: frame_threads_0222 (RW)
0xdf: frame_threads_0223 (RW)
0xe0: frame_threads_0224 (RW)
0xe1: frame_threads_0225 (RW)
0xe2: frame_threads_0226 (RW)
0xe3: frame_threads_0227 (RW)
0xe4: frame_threads_0228 (RW)
0xe5: frame_threads_0229 (RW)
0xe6: frame_threads_0230 (RW)
0xe7: frame_threads_0231 (RW)
0xe8: frame_threads_0232 (RW)
0xe9: frame_threads_0233 (RW)
0xea: frame_threads_0234 (RW)
0xeb: frame_threads_0235 (RW)
0xec: frame_threads_0236 (RW)
0xed: frame_threads_0237 (RW)
0xee: frame_threads_0238 (RW)
0xef: frame_threads_0239 (RW)
0xf0: frame_threads_0240 (RW)
0xf1: frame_threads_0241 (RW)
0xf2: frame_threads_0242 (RW)
0xf3: frame_threads_0243 (RW)
0xf4: frame_threads_0244 (RW)
0xf5: frame_threads_0245 (RW)
0xf6: frame_threads_0246 (RW)
0xf7: frame_threads_0247 (RW)
0xf8: frame_threads_0248 (RW)
0xf9: frame_threads_0249 (RW)
0xfa: frame_threads_0250 (RW)
0xfb: frame_threads_0251 (RW)
0xfc: frame_threads_0252 (RW)
0xfd: frame_threads_0253 (RW)
0xfe: frame_threads_0254 (RW)
0xff: frame_threads_0255 (RW)
0x100: frame_threads_0256 (RW)
0x101: frame_threads_0257 (RW)
0x102: frame_threads_0258 (RW)
0x103: frame_threads_0259 (RW)
0x104: frame_threads_0260 (RW)
0x105: frame_threads_0261 (RW)
0x106: frame_threads_0262 (RW)
0x107: frame_threads_0263 (RW)
0x108: frame_threads_0264 (RW)
0x109: frame_threads_0265 (RW)
0x10a: frame_threads_0266 (RW)
0x10b: frame_threads_0267 (RW)
0x10c: frame_threads_0268 (RW)
0x10d: frame_threads_0269 (RW)
0x10e: frame_threads_0270 (RW)
0x10f: frame_threads_0271 (RW)
0x110: frame_threads_0272 (RW)
0x111: frame_threads_0273 (RW)
0x112: frame_threads_0274 (RW)
0x113: frame_threads_0275 (RW)
0x114: frame_threads_0276 (RW)
0x115: frame_threads_0277 (RW)
0x116: frame_threads_0278 (RW)
0x117: frame_threads_0279 (RW)
0x118: frame_threads_0280 (RW)
0x119: frame_threads_0281 (RW)
0x11a: frame_threads_0282 (RW)
0x11b: frame_threads_0283 (RW)
0x11c: frame_threads_0284 (RW)
0x11d: frame_threads_0285 (RW)
0x11e: frame_threads_0286 (RW)
0x11f: frame_threads_0287 (RW)
0x120: frame_threads_0288 (RW)
0x121: frame_threads_0289 (RW)
0x122: frame_threads_0290 (RW)
0x123: frame_threads_0291 (RW)
0x124: frame_threads_0292 (RW)
0x125: frame_threads_0293 (RW)
0x126: frame_threads_0294 (RW)
0x127: frame_threads_0295 (RW)
0x128: frame_threads_0296 (RW)
0x129: frame_threads_0297 (RW)
0x12a: frame_threads_0298 (RW)
0x12b: frame_threads_0299 (RW)
0x12c: frame_threads_0300 (RW)
0x12d: frame_threads_0301 (RW)
0x12e: frame_threads_0302 (RW)
0x12f: frame_threads_0303 (RW)
0x130: frame_threads_0304 (RW)
0x131: frame_threads_0305 (RW)
0x132: frame_threads_0306 (RW)
0x133: frame_threads_0307 (RW)
0x134: frame_threads_0308 (RW)
0x135: frame_threads_0309 (RW)
0x136: frame_threads_0310 (RW)
0x137: frame_threads_0311 (RW)
0x138: frame_threads_0312 (RW)
0x139: frame_threads_0313 (RW)
0x13a: frame_threads_0314 (RW)
0x13b: frame_threads_0315 (RW)
0x13c: frame_threads_0316 (RW)
0x13d: frame_threads_0317 (RW)
0x13e: frame_threads_0318 (RW)
0x13f: frame_threads_0319 (RW)
0x140: frame_threads_0320 (RW)
0x141: frame_threads_0321 (RW)
0x142: frame_threads_0322 (RW)
0x143: frame_threads_0323 (RW)
0x144: frame_threads_0324 (RW)
}
tcb_threads {
cspace: cnode_threads (guard: 0, guard_size: 60)
ipc_buffer_slot: ipc_threads_obj (RW)
vspace: vspace_threads
}
vspace_threads {
0x0: pdpt_threads_0000
}
}

irq maps {

}